###############################################################################
#TSMC Library/IP Product
#Filename: antenna_8.lef
#Technology: CL013G
#Product Type: Standard I/O
#Product Name: tpd013n3
#Version: 210a
###############################################################################
# 
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
# 
###############################################################################

jjfwjfwjjfwjfwjjfwjfwjjfwjfwjjfwjfwjjfwjfwjjfwjfwjjfwjfwjjfwjfwjjfwjfw